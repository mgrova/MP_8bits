-- This behavior can be modeled using an RTL process that uses the address bus and the 
-- write signal to create a synchronous enable condition. 
-- Each port is modeled with its own process. The following VHDL shows how the output ports at

